module page_sexa_bb(
    input wire clk_0,
    input wire [48 : 0] din_leaf_bft2interface_0,
    output wire  [48 : 0] dout_leaf_interface2bft_0,
    input wire resend_0,
    input wire reset_0,
    input wire ap_start_0,

    input wire clk_1,
    input wire [48 : 0] din_leaf_bft2interface_1,
    output wire  [48 : 0] dout_leaf_interface2bft_1,
    input wire resend_1,
    input wire reset_1,
    input wire ap_start_1,

    input wire clk_2,
    input wire [48 : 0] din_leaf_bft2interface_2,
    output wire  [48 : 0] dout_leaf_interface2bft_2,
    input wire resend_2,
    input wire reset_2,
    input wire ap_start_2,

    input wire clk_3,
    input wire [48 : 0] din_leaf_bft2interface_3,
    output wire  [48 : 0] dout_leaf_interface2bft_3,
    input wire resend_3,
    input wire reset_3,
    input wire ap_start_3,

    input wire clk_4,
    input wire [48 : 0] din_leaf_bft2interface_4,
    output wire  [48 : 0] dout_leaf_interface2bft_4,
    input wire resend_4,
    input wire reset_4,
    input wire ap_start_4,

    input wire clk_5,
    input wire [48 : 0] din_leaf_bft2interface_5,
    output wire  [48 : 0] dout_leaf_interface2bft_5,
    input wire resend_5,
    input wire reset_5,
    input wire ap_start_5
    );
   
endmodule
